module Ahbmli(
    output[7:0] io_out
);



  assign io_out = 8'h2a;
endmodule

